.PS
cct_init
resistor(down_)
.PE

